LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;
ENTITY InstructionM_E IS
PORT (
address : IN std_logic_vector(31 downto 0);
dataout : OUT std_logic_vector(31 downto 0)
);
END ENTITY InstructionM_E;

ARCHITECTURE InstructionM_A OF InstructionM_E IS 
TYPE ram_type IS ARRAY(0 TO 75) of std_logic_vector(15 DOWNTO 0);
SIGNAL RAM : ram_type:=(
--std_logic_vector(to_unsigned(0,16)), std_logic_vector(to_unsigned(1,16)), std_logic_vector(to_unsigned(2,16)), 
--std_logic_vector(to_unsigned(3,16)), std_logic_vector(to_unsigned(4,16)), std_logic_vector(to_unsigned(5,16))

"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0101010111110010",
"0101010111110011",
"0101010111110100",
"1110010011110001",
"0000000000000101",

"0000000000000000",	-- NOP
"0000000000000000",	-- NOP

"0010001011110001",
"0010001011110010",
"0010001111110001",
"0010001111110010",
"0101010111110101",

"0000000000000000",	-- NOP
"0000000000000000",	-- NOP

"1110111001010010",
"0000000011001000",
"1110111001010001",
"0000000011001010",
"1110110101010011",
"0000000011001010",
"1110110101010100",
"0000000011001000",



"0000000000000000",	-- NOP

------------------------------


"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000"	-- NOP

);
BEGIN
	dataout <= RAM(to_integer(unsigned(address(18 downto 0))))& RAM(to_integer(unsigned(address(18 downto 0)))+1);
			
END InstructionM_A;