LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;
ENTITY InstructionM_E IS
PORT (
address : IN std_logic_vector(31 downto 0);
dataout : OUT std_logic_vector(31 downto 0)
);
END ENTITY InstructionM_E;

ARCHITECTURE InstructionM_A OF InstructionM_E IS 
TYPE ram_type IS ARRAY(0 TO 61) of std_logic_vector(15 DOWNTO 0);
SIGNAL RAM : ram_type:=(
--std_logic_vector(to_unsigned(0,16)), std_logic_vector(to_unsigned(1,16)), std_logic_vector(to_unsigned(2,16)), 
--std_logic_vector(to_unsigned(3,16)), std_logic_vector(to_unsigned(4,16)), std_logic_vector(to_unsigned(5,16))

"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",

"0101010111110010", -- IN R2

"0000000000000000",
"0000000000000000",

"1001011000100010",	-- SHL R2,2
"0000000010000000",

"0000000000000000",	-- NOP
"0000000000000000",	-- NOP

"1001011100100010", -- SHR R2,3
"0000000011000000",

"0000000000000000",	-- NOP
"0000000000000000",	-- NOP

"1110011100100010", -- IADD R2, FFFF
"1111111111111111",

"0000000000000000",	-- NOP
"0000000000000000",	-- NOP

"1110010000010001", -- LDM r1, 1
"0000000000000001",

"0001111100010010", -- ADD R1,R2



"0000000000000000",	-- NOP

------------------------------

"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000",	-- NOP
"0000000000000000"	-- NOP

);
BEGIN
	dataout <= RAM(to_integer(unsigned(address(18 downto 0))))& RAM(to_integer(unsigned(address(18 downto 0)))+1);
			
END InstructionM_A;